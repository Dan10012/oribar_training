
package functions;

	function byte[16] sub_bytes_func (byte[16] state_data);

	endfunction 

endpackage